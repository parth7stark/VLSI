`include "sixtyfourBitAdder.v"

module top;
	reg[63:0] A,B;
	reg Cin;
	wire[63:0] sum;
	wire Cout;
	
	sixtyfourBitAdder F0(A,B,Cin,sum,Cout);
	
	initial 
	begin
		
		A= {$random}%(2**64-1);
		B= {$random}%(10000);
		Cin =0;
		#10
		A = 64'b0000000000000000000000000000000000000000000000000000000000000000 ; B = 64'b0000000000000000000000000000000000000000000000000000000000000000; Cin = 0;
		
		#10 A = 64'b0011000000000000000000000000000000000000000000000000000000000000; B = 64'b0100000000000000000000000000000000000000000000000000000000000000;
		#10 A = 64'b0111101000010100000000000000000011111111111111111111111111111111; B = 64'b0110011000000110000000000000000011111111111111111111111111111111; Cin = 1;
		#10 A = 64'b1111111111111111111111111111111111111111111111111111111111111111; B = 64'b1111111111111111111111111111111111111111111111111111111111111111;
	end
	
	
	
	initial
	begin
		$monitor($time, " A = %d, B = %d, Cin = %d, Sum = %d, ca = %d",A,B,Cin,sum, Cout);
		$dumpfile("64BitAdder.vcd");
		$dumpvars;
	end

endmodule	
